module AsyncFIFO (
    input wire clk_write,
    input wire clk_read,
    input wire rst,
    input wire [7:0] data_in,
    input wire write_enable,
    input wire read_enable,
    output logic [7:0] data_out,
    output logic full,
    output logic empty,
    output logic almost_full,
    output logic almost_empty
):



endmodule

