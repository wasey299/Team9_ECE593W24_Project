import uvm_pkg::*;
`include "uvm_macros.svh"
`include "fifo_if.sv"
`include "trans.sv"
`include "w_trans.sv"
`include "wr_config.sv"
`include "rd_config.sv"
`include "env_config.sv"
`include "wr_driver.sv"
`include "wr_monitor.sv"
`include "wr_sequencer.sv"
`include "wr_agent.sv"
`include "w_sequence.sv"
`include "rd_driver.sv"
`include "rd_monitor.sv"
`include "rd_sequencer.sv"
`include "rd_agent.sv"
`include "r_sequence.sv"
`include "v_sequencer.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "v_sequence.sv"
`include "test.sv"
`include "top.sv"