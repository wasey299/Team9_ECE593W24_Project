module AsyncFIFO (
    input wire clk_write,
    input wire clk_read,
    input wire rst,
    input wire [7:0] data_in,
    input wire write_enable,
    input wire read_enable,
    output logic [7:0] data_out,
    output logic full,
    output logic empty,
    output logic almost_full,
    output logic almost_empty
):

parameter DEPTH = 256; 

reg [7:0] memory [0:DEPTH-1];
reg [$clog2(DEPTH):0] front_index, rear_index;
reg [$clog2(DEPTH):0] next_rear_index;
reg [$clog2(DEPTH):0] count;










endmodule

